`timescale 1ns / 1ps

module comparator_32_bit (
  input [31:0] A,
  input [31:0] B,
  output EQ,
  output GT,
  output LT
);

wire [31:0] xor_result;

assign xor_result = A ^ B;

// Calculate equality
assign EQ = ~(|xor_result);

// Calculate greater than (GT) - Explicitly define outputs for all bits
wire GT_0, GT_1, GT_2, GT_3, GT_4, GT_5, GT_6, GT_7,
    GT_8, GT_9, GT_10, GT_11, GT_12, GT_13, GT_14, GT_15, 
    GT_16, GT_17, GT_18, GT_19, GT_20, GT_21, GT_22, GT_23, 
    GT_24, GT_25, GT_26, GT_27, GT_28, GT_29, GT_30, GT_31;
    
  // Compare MSB (Most Significant Bit)
assign GT_31 = (~A[31] & B[31]);

// Compare remaining bits (30 to 0)
assign GT_30 = ~A[31] & (A[30] ^ B[30]);
assign GT_29 = (~A[31] & ~A[30]) & (A[29] ^ B[29]);
assign GT_28 = (~A[31] & ~A[30] & ~A[29]) & (A[28] ^ B[28]);
assign GT_27 = (~A[31] & ~A[30] & ~A[29] & ~A[28]) & (A[27] ^ B[27]);
assign GT_26 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27]) & (A[26] ^ B[26]);
assign GT_25 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26]) & (A[25] ^ B[25]);
assign GT_24 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25]) & (A[24] ^ B[24]);
assign GT_23 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24]) & (A[23] ^ B[23]);
assign GT_22 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23]) & (A[22] ^ B[22]);
assign GT_21 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22]) & (A[21] ^ B[21]);
assign GT_20 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21]) & (A[20] ^ B[20]);
assign GT_19 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20]) & (A[19] ^ B[19]);
assign GT_18 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19]) & (A[18] ^ B[18]);
assign GT_17 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18]) & (A[17] ^ B[17]);
assign GT_16 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17]) & (A[16] ^ B[16]);
assign GT_15 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16]) & (A[15] ^ B[15]);
assign GT_14 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15]) & (A[14] ^ B[14]);
assign GT_13 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14]) & (A[13] ^ B[13]);
assign GT_12 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13]) & (A[12] ^ B[12]);
assign GT_11 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12]) & (A[11] ^ B[11]);
assign GT_10 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11]) & (A[10] ^ B[10]);
assign GT_9 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10]) & (A[9] ^ B[9]);
assign GT_8 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9]) & (A[8] ^ B[8]);
assign GT_7 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8]) & (A[7] ^ B[7]);
assign GT_6 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7]) & (A[6] ^ B[6]);
assign GT_5 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6]) & (A[5] ^ B[5]);
assign GT_4 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5]) & (A[4] ^ B[4]);
assign GT_3 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4]) & (A[3] ^ B[3]);
assign GT_2 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3]) & (A[2] ^ B[2]);
assign GT_1 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & ~A[2]) & (A[1] ^ B[1]);
assign GT_0 = (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & ~A[2] & ~A[1]) & (A[0] ^ B[0]);

// Assign GT output based on individual bit comparisons
  assign GT = GT_0 | GT_1 | GT_2 | GT_3 | GT_4 | GT_5 | GT_6 | GT_7 |
              GT_8 | GT_9 | GT_10 | GT_11 | GT_12 | GT_13 | GT_14 | 
              GT_15 | GT_16 | GT_17 | GT_18 | GT_19 | GT_20 | GT_21 |
              GT_22 | GT_23 | GT_24 | GT_25 | GT_26 | GT_27 | GT_28 |
              GT_29 | GT_30 | GT_31;
              
// Calculate less than (LT) - Similar logic as GT, but using opposite logic for A and B
wire LT_0, LT_1, LT_2, LT_3, LT_4, LT_5, LT_6, LT_7,
     LT_8, LT_9, LT_10, LT_11, LT_12, LT_13, LT_14, LT_15,
     LT_16, LT_17, LT_18, LT_19, LT_20, LT_21, LT_22, LT_23,
     LT_24, LT_25, LT_26, LT_27, LT_28, LT_29, LT_30, LT_31;
     
// Compare MSB
assign LT_31 = (A[31] & ~B[31]);

// Compare remaining bits
assign LT_30 = (A[31] & ~A[30] & B[30]) | (~A[31] & ~B[31] & (A[30] ^ B[30]));
assign LT_29 = (A[31] & ~A[30] & ~A[29] & B[29]) | (~A[31] & ~A[30] & ~B[30] & (A[29] ^ B[29]));
assign LT_28 = (A[31] & ~A[30] & ~A[29] & ~A[28] & B[28]) | (~A[31] & ~A[30] & ~A[29] & ~B[29] & (A[28] ^ B[28]));
assign LT_27 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & B[27]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~B[28] & (A[27] ^ B[27]));
assign LT_26 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & B[26]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~B[27] & (A[26] ^ B[26]));
assign LT_25 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & B[25]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~B[26] & (A[25] ^ B[25]));
assign LT_24 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & B[24]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~B[25] & (A[24] ^ B[24]));
assign LT_23 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & B[23]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~B[24] & (A[23] ^ B[23]));
assign LT_22 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & B[22]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~B[23] & (A[22] ^ B[22]));
assign LT_21 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & B[21]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~B[22] & (A[21] ^ B[21]));
assign LT_20 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & B[20]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~B[21] & (A[20] ^ B[20]));
assign LT_19 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & B[19]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~B[20] & (A[19] ^ B[19]));
assign LT_18 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & B[18]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~B[19] & (A[18] ^ B[18]));
assign LT_17 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & B[17]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~B[18] & (A[17] ^ B[17]));
assign LT_16 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & B[16]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[16] ^ B[16]));
assign LT_15 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & B[16]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[16] ^ B[16]));
assign LT_14 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & B[15]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[15] ^ B[15]));
assign LT_13 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & B[14]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[14] ^ B[14]));
assign LT_12 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & B[13]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[13] ^ B[13]));
assign LT_11 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & B[12]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[12] ^ B[12]));
assign LT_10 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & B[11]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[11] ^ B[11]));
assign LT_9 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & B[10]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[10] ^ B[10]));
assign LT_8 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & B[9]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[9] ^ B[9]));
assign LT_7 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & B[8]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[8] ^ B[8]));
assign LT_6 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & B[7]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[7] ^ B[7]));
assign LT_5 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & B[6]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[6] ^ B[6]));
assign LT_4 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & B[5]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[5] ^ B[5]));
assign LT_3 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & B[4]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[4] ^ B[4]));
assign LT_2 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & B[3]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[3] ^ B[3]));
assign LT_1 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & ~A[2] & B[2]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[2] ^ B[2]));
assign LT_0 = (A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & ~A[2] & ~A[1] & B[1]) | (~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~B[17] & (A[1] ^ B[1]));

 // Assign LT output based on individual bit comparisons
  assign LT = LT_0 | LT_1 | LT_2 | LT_3 | LT_4 | LT_5 | LT_6 | LT_7 |
              LT_8 | LT_9 | LT_10 | LT_11 | LT_12 | LT_13 | LT_14 | LT_15 |
              LT_16 | LT_17 | LT_18 | LT_19 | LT_20 | LT_21 | LT_22 | LT_23 | 
              LT_24 | LT_25 | LT_26 | LT_27 | LT_28 | LT_29 | LT_30 | LT_31;

endmodule

