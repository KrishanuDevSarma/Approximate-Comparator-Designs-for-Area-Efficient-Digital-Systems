`timescale 1ns / 1ps

module approx_comparator_32_bit (
  input [31:0] A,
  input [31:0] B,
  output EQ,
  output reg GT,
  output reg LT
);

  wire [31:0] xor_result;

  // Calculate XOR of A and B
  assign xor_result = A ^ B;

  // Calculate equality
  assign EQ = |(xor_result);

  // Calculate greater than (GT)
  always @* begin
    GT = &(~A[31] & B[31]) | (~A[31] & (A[30] ^ B[30])) | ((~A[31] & ~A[30]) & (A[29] ^ B[29])) | 
     (((~A[31] & ~A[30] & ~A[29]) & (A[28] ^ B[28]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28]) & (A[27] ^ B[27]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27]) & (A[26] ^ B[26]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26]) & (A[25] ^ B[25]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25]) & (A[24] ^ B[24]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24]) & (A[23] ^ B[23]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23]) & (A[22] ^ B[22]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22]) & (A[21] ^ B[21]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21]) & (A[20] ^ B[20]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20]) & (A[19] ^ B[19]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19]) & (A[18] ^ B[18]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18]) & (A[17] ^ B[17]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17]) & (A[16] ^ B[16]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16]) & (A[15] ^ B[15]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15]) & (A[14] ^ B[14]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14]) & (A[13] ^ B[13]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13]) & (A[12] ^ B[12]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12]) & (A[11] ^ B[11]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11]) & (A[10] ^ B[10]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10]) & (A[9] ^ B[9]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9]) & (A[8] ^ B[8]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8]) & (A[7] ^ B[7]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7]) & (A[6] ^ B[6]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6]) & (A[5] ^ B[5]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5]) & (A[4] ^ B[4]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4]) & (A[3] ^ B[3]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3]) & (A[2] ^ B[2]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & ~A[2]) & (A[1] ^ B[1]))) |
     (((~A[31] & ~A[30] & ~A[29] & ~A[28] & ~A[27] & ~A[26] & ~A[25] & ~A[24] & ~A[23] & ~A[22] & ~A[21] & ~A[20] & ~A[19] & ~A[18] & ~A[17] & ~A[16] & ~A[15] & ~A[14] & ~A[13] & ~A[12] & ~A[11] & ~A[10] & ~A[9] & ~A[8] & ~A[7] & ~A[6] & ~A[5] & ~A[4] & ~A[3] & ~A[2] & ~A[1]) & (A[0] ^ B[0])));
 // Continue pattern for all 32 bits
  end

  // Calculate less than (LT)
  always @* begin
    LT = ((A[31] & ~B[31]) |
      (A[31] & (~A[30] ^ B[30])) |
      ((A[31] & A[30]) & (~A[29] ^ B[29])) |
      ((A[31] & A[30] & A[29]) & (~A[28] ^ B[28])) |
      ((A[31] & A[30] & A[29] & A[28]) & (~A[27] ^ B[27])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27]) & (~A[26] ^ B[26])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26]) & (~A[25] ^ B[25])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25]) & (~A[24] ^ B[24])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24]) & (~A[23] ^ B[23])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23]) & (~A[22] ^ B[22])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22]) & (~A[21] ^ B[21])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21]) & (~A[20] ^ B[20])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20]) & (~A[19] ^ B[19])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19]) & (~A[18] ^ B[18])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18]) & (~A[17] ^ B[17])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17]) & (~A[16] ^ B[16])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16]) & (~A[15] ^ B[15])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15]) & (~A[14] ^ B[14])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14]) & (~A[13] ^ B[13])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13]) & (~A[12] ^ B[12])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12]) & (~A[11] ^ B[11])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11]) & (~A[10] ^ B[10])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10]) & (~A[9] ^ B[9])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9]) & (~A[8] ^ B[8])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8]) & (~A[7] ^ B[7])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7]) & (~A[6] ^ B[6])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7] & A[6]) & (~A[5] ^ B[5])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7] & A[6] & A[5]) & (~A[4] ^ B[4])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7] & A[6] & A[5] & A[4]) & (~A[3] ^ B[3])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7] & A[6] & A[5] & A[4] & A[3]) & (~A[2] ^ B[2])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7] & A[6] & A[5] & A[4] & A[3] & A[2]) & (~A[1] ^ B[1])) |
      ((A[31] & A[30] & A[29] & A[28] & A[27] & A[26] & A[25] & A[24] & A[23] & A[22] & A[21] & A[20] & A[19] & A[18] & A[17] & A[16] & A[15] & A[14] & A[13] & A[12] & A[11] & A[10] & A[9] & A[8] & A[7] & A[6] & A[5] & A[4] & A[3] & A[2] & A[1]) & (~A[0] ^ B[0])) |
      1'b0);
// Continue pattern for all 32 bits
  end

endmodule
